`include "main.v"

module main_tb();
    
endmodule